`default_nettype none

module Clock(
  output logic clock,
  input logic halt
);

endmodule